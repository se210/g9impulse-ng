sdram_pll_inst : sdram_pll PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig,
		c1	 => c1_sig,
		locked	 => locked_sig
	);
